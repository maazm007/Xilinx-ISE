module not_gate(x,out);
	input x;
	output out;
	assign out = ~x;
endmodule
